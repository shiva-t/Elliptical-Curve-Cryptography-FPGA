module inverse(out,a,f,clock);
output reg [3:0]out;
input [3:0]a;
input [4:0]f;
input clock;

reg [3:0]u;
reg [4:0]v;
reg [4:0]g1=5'd1;
reg [4:0]g2=5'd0;
//reg begin_s=1;

always@(a)
begin
u=a; v=f;
g1=5'd1;g2=5'd0;
end 

always@(posedge clock)
begin 

if ( (u[3]==1) | (u[2]==1) | (u[1]==1) | (v[4]==1) | (v[3]==1) | (v[2]==1) | (v[1]==1)  )   //While (u!=1and v!=1)
begin

	if(u[0]==0 & ((u[3]==1) | (u[2]==1) | (u[1]==1)))   //3.1
	begin
		u[0]=u[1];
		u[1]=u[2];
		u[2]=u[3];
		u[3]=1'b0;

		if(g1[0]==0 & ( (g1[1]==1) | (g1[2]==1) | (g1[3]==1) | (g1[4]==1) ) )

		begin
			g1[0]=g1[1];   //divide by z
			g1[1]=g1[2];
			g1[2]=g1[3];
			g1[3]=g1[4];
			g1[4]=1'b0;


		end
		else 
		begin
			

			g1[0]=g1[0]^ f[0];
			g1[1]=g1[1]^ f[1];
			g1[2]=g1[2]^ f[2];
			g1[3]=g1[3]^ f[3];
			g1[4]=g1[4]^ f[4];

			

			g1[0]=g1[1];   //divide by z
			g1[1]=g1[2];
			g1[2]=g1[3];
			g1[3]=g1[4];
			g1[4]=1'b0;
		end
	end     //end of 3.1

	if(u[0]==0 & ((u[3]==1) | (u[2]==1) | (u[1]==1)))   //3.1
	begin
		u[0]=u[1];
		u[1]=u[2];
		u[2]=u[3];
		u[3]=1'b0;

		if(g1[0]==0 & ( (g1[1]==1) | (g1[2]==1) | (g1[3]==1) | (g1[4]==1) ) )

		begin
			g1[0]=g1[1];   //divide by z
			g1[1]=g1[2];
			g1[2]=g1[3];
			g1[3]=g1[4];
			g1[4]=1'b0;


		end
		else 
		begin
			
			g1[0]=g1[0]^ f[0];
			g1[1]=g1[1]^ f[1];
			g1[2]=g1[2]^ f[2];
			g1[3]=g1[3]^ f[3];
			g1[4]=g1[4]^ f[4];


			g1[0]=g1[1];   //divide by z
			g1[1]=g1[2];
			g1[2]=g1[3];
			g1[3]=g1[4];
			g1[4]=1'b0;
		end
	end  

	if(u[0]==0 & ((u[3]==1) | (u[2]==1) | (u[1]==1)))   //3.1
	begin
		u[0]=u[1];
		u[1]=u[2];
		u[2]=u[3];
		u[3]=1'b0;

		if(g1[0]==0 & ( (g1[1]==1) | (g1[2]==1) | (g1[3]==1) | (g1[4]==1) ) )

		begin
			g1[0]=g1[1];   //divide by z
			g1[1]=g1[2];
			g1[2]=g1[3];
			g1[3]=g1[4];
			g1[4]=1'b0;


		end
		else 
		begin
			
			g1[0]=g1[0]^ f[0];
			g1[1]=g1[1]^ f[1];
			g1[2]=g1[2]^ f[2];
			g1[3]=g1[3]^ f[3];
			g1[4]=g1[4]^ f[4];


			g1[0]=g1[1];   //divide by z
			g1[1]=g1[2];
			g1[2]=g1[3];
			g1[3]=g1[4];
			g1[4]=1'b0;
		end
	end  

	
	if(v[0]==0 & ((v[4]==1) | (v[3]==1) | (v[2]==1) | (v[1]==1)))   //3.2
	begin
		v[0]=v[1];
		v[1]=v[2];
		v[2]=v[3];
		v[3]=v[4];
		v[4]=1'b0;

		if(g2[0]==0 & ( (g2[1]==1) | (g2[2]==1) | (g2[3]==1) | (g2[4]==1) ) )

		begin
			g2[0]=g2[1];   //divide by z
			g2[1]=g2[2];
			g2[2]=g2[3];
			g2[3]=g2[4];
			g2[4]=1'b0;


		end
		else 
		begin
			
			g2[0]=g2[0]^ f[0];
			g2[1]=g2[1]^ f[1];
			g2[2]=g2[2]^ f[2];
			g2[3]=g2[3]^ f[3];
			g2[4]=g2[4]^ f[4];


			g2[0]=g2[1];   //divide by z
			g2[1]=g2[2];
			g2[2]=g2[3];
			g2[3]=g2[4];
			g2[4]=1'b0;
		end
	end     //end of 3.2

	if(v[0]==0 & ((v[4]==1) | (v[3]==1) | (v[2]==1) | (v[1]==1)))   //3.2
	begin
		v[0]=v[1];
		v[1]=v[2];
		v[2]=v[3];
		v[3]=v[4];
		v[4]=1'b0;

		if(g2[0]==0 & ( (g2[1]==1) | (g2[2]==1) | (g2[3]==1) | (g2[4]==1) ) )

		begin
			g2[0]=g2[1];   //divide by z
			g2[1]=g2[2];
			g2[2]=g2[3];
			g2[3]=g2[4];
			g2[4]=1'b0;


		end
		else 
		begin
			
			g2[0]=g2[0]^ f[0];
			g2[1]=g2[1]^ f[1];
			g2[2]=g2[2]^ f[2];
			g2[3]=g2[3]^ f[3];
			g2[4]=g2[4]^ f[4];

			g2[0]=g2[1];   //divide by z
			g2[1]=g2[2];
			g2[2]=g2[3];
			g2[3]=g2[4];
			g2[4]=1'b0;
		end
	end     //end of 3.2

	if(v[0]==0 & ((v[4]==1) | (v[3]==1) | (v[2]==1) | (v[1]==1)))   //3.2
	begin
		v[0]=v[1];
		v[1]=v[2];
		v[2]=v[3];
		v[3]=v[4];
		v[4]=1'b0;

		if(g2[0]==0 & ( (g2[1]==1) | (g2[2]==1) | (g2[3]==1) | (g2[4]==1) ) )

		begin
			g2[0]=g2[1];   //divide by z
			g2[1]=g2[2];
			g2[2]=g2[3];
			g2[3]=g2[4];
			g2[4]=1'b0;


		end
		else 
		begin
			
			g2[0]=g2[0]^ f[0];
			g2[1]=g2[1]^ f[1];
			g2[2]=g2[2]^ f[2];
			g2[3]=g2[3]^ f[3];
			g2[4]=g2[4]^ f[4];

			g2[0]=g2[1];   //divide by z
			g2[1]=g2[2];
			g2[2]=g2[3];
			g2[3]=g2[4];
			g2[4]=1'b0;
		end
	end     //end of 3.2

	//3.3
	if( ((u[3]==1) & (v[4]==0) & (v[3]==0)) | ( (u[3]==0) & (u[2]==1) & (v[4]==0) & (v[3]==0) & (v[2]==0)) | ( (u[3]==0) & (u[2]==0) & (u[1]==1) & (v[4]==0) & (v[3]==0) & (v[2]==0) & (v[1]==0))  |   
	( (u[3]==0) & (u[2]==0) & (u[1]==0) & (u[0]==1) & (v[4]==0) & (v[3]==0) & (v[2]==0) & (v[1]==0) & (v[0]==0))     )
	begin

		u[0]=u[0]^ v[0];
		u[1]=u[1]^ v[1];
		u[2]=u[2]^ v[2];
		u[3]=u[3]^ v[3];
		

		g1[0]=g2[0]^ g1[0];
		g1[1]=g2[1]^ g1[1];
		g1[2]=g2[2]^ g1[2];
		g1[3]=g2[3]^ g1[3];
		g1[4]=g2[4]^ g1[4];	

	end
	else begin
		
		v[0]=v[0] ^ u[0];
		v[1]=v[1] ^ u[1];
		v[2]=v[2] ^ u[2];
		v[3]=v[3] ^ u[3];		
		
		g2[0]=g2[0]^ g1[0];
		g2[1]=g2[1]^ g1[1];
		g2[2]=g2[2]^ g1[2];
		g2[3]=g2[3]^ g1[3];
		g2[4]=g2[4]^ g1[4];

	end //3.3 ends

	//if((u[3]==0) & (u[2]==0) & (u[1]==0) & (v[3]==0) & (v[2]==0) & (v[1]==0) & (v[4]==0)  )
	if( ((u==4'b0001) & (v==5'b00000)) | ((u==4'b0000) & (v==5'b00001)) )begin
	if(u==4'b0001)
	begin
		out=g1;
	end
	else out=g2;
	end

end


end

endmodule 


module tb_inverse();
wire [3:0]out;
reg [3:0]a;
reg [4:0]f;
reg clock;
inverse uut(.out(out),.a(a),.f(f),.clock(clock));
initial forever #5 clock=~clock;

initial begin
//clock=1'b0;a=4'b0100; f=5'b10011;
//clock=1'b0;a=4'b1001; f=5'b10011;
//clock=1'b0;a=4'b1001; f=5'b10011;
clock=1'b1;a=4'b1111; f=5'b10011;
//#50 a=4'b1001;
#300 $stop;
end


endmodule 